��  CCircuit��  CSerializeHack           ��  CPart              ���  CMotorEM�� 	 CTerminal  `�a�                �          
�  `�a�                           �� 	 CMechTerm       �                                  l�q�     	        �            T�l�         ��      bK�6�>       �                       �        ��  CSPST��  CToggle   � �         
�  � ��             "@          
�  �1�               �            ��           ��    ��  CBattery��  CValue  � �� �    9V(          "@      �? V 
�  � �� �              "@          
�  � �� �                            � �� �         ��                    ���  CWire  � �a�       �  0�a�      �  � �� �                    �                                                                  �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 